// systolic_top.v
// Top-level: classic 2D systolic array + small controller.
// Expects A (ROWS x K) and B (K x COLS) as flattened int8 matrices.
// Produces C (ROWS x COLS) as flattened int32 matrix.

module systolic_top #(
    parameter DATA_W = 8,
    parameter ACC_W  = 32,
    parameter ROWS   = 4,
    parameter COLS   = 4,
    parameter K      = 4
)(
    input  wire clk,
    input  wire rst_n,

    input  wire start,
    output wire busy,
    output wire done,

    input  wire signed [ROWS*K*DATA_W-1:0] a_flat,
    input  wire signed [K*COLS*DATA_W-1:0] b_flat,

    output reg  signed [ROWS*COLS*ACC_W-1:0] c_flat
);

    // internal storage for A and B
    integer r, c;

    reg signed [DATA_W-1:0] A_reg [0:ROWS-1][0:K-1];
    reg signed [DATA_W-1:0] B_reg [0:K-1][0:COLS-1];

    // controller
    wire ctrl_busy;
    wire ctrl_done;
    wire valid_src;
    wire [$clog2(K):0] k_idx;

    systolic_controller #(
        .ROWS(ROWS),
        .COLS(COLS),
        .K   (K)
    ) u_ctrl (
        .clk      (clk),
        .rst_n    (rst_n),
        .start    (start),
        .busy     (ctrl_busy),
        .done     (ctrl_done),
        .valid_src(valid_src),
        .k_idx    (k_idx)
    );

    assign busy = ctrl_busy;
    assign done = ctrl_done;

    // build A/B input buses for systolic_array
    reg signed [ROWS*DATA_W-1:0] a_in_bus;
    reg signed [COLS*DATA_W-1:0] b_in_bus;

    // outputs from array
    wire signed [ROWS*COLS*ACC_W-1:0] c_bus;
    wire [ROWS*COLS-1:0]              c_valid;

    systolic_array #(
        .DATA_W(DATA_W),
        .ACC_W (ACC_W),
        .ROWS  (ROWS),
        .COLS  (COLS)
    ) u_array (
        .clk     (clk),
        .rst_n   (rst_n),
        .valid_in(valid_src),
        .a_in_bus(a_in_bus),
        .b_in_bus(b_in_bus),
        .c_bus   (c_bus),
        .c_valid (c_valid)
    );

    // flags to capture each C(i,j) only once
    reg [ROWS*COLS-1:0] captured;

    // unpack A_flat and B_flat once when we get a start pulse in IDLE
    // here, we simply load every time start is seen while not busy
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for (r = 0; r < ROWS; r = r + 1) begin
                for (c = 0; c < K; c = c + 1) begin
                    A_reg[r][c] <= '0;
                end
            end
            for (r = 0; r < K; r = r + 1) begin
                for (c = 0; c < COLS; c = c + 1) begin
                    B_reg[r][c] <= '0;
                end
            end
        end else begin
            if (start && !ctrl_busy) begin
                // load A
                for (r = 0; r < ROWS; r = r + 1) begin
                    for (c = 0; c < K; c = c + 1) begin
                        int idx;
                        idx = r*K + c;
                        A_reg[r][c] <= a_flat[(idx+1)*DATA_W-1 -: DATA_W];
                    end
                end

                // load B
                for (r = 0; r < K; r = r + 1) begin
                    for (c = 0; c < COLS; c = c + 1) begin
                        int idx;
                        idx = r*COLS + c;
                        B_reg[r][c] <= b_flat[(idx+1)*DATA_W-1 -: DATA_W];
                    end
                end

                // reset capture flags and C outputs
                captured <= '0;
                c_flat   <= '0;
            end
        end
    end

    // drive left and top edge inputs to systolic_array
    always @(*) begin
        a_in_bus = '0;
        b_in_bus = '0;

        if (ctrl_busy && (k_idx < K)) begin
            // use k_idx as the column index in A, row index in B
            for (r = 0; r < ROWS; r = r + 1) begin
                a_in_bus[(r+1)*DATA_W-1 -: DATA_W] = A_reg[r][k_idx];
            end
            for (c = 0; c < COLS; c = c + 1) begin
                b_in_bus[(c+1)*DATA_W-1 -: DATA_W] = B_reg[k_idx][c];
            end
        end
    end

    // capture C outputs when each PE asserts its valid for the first time
    integer idx;
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            captured <= '0;
            c_flat   <= '0;
        end else begin
            for (idx = 0; idx < ROWS*COLS; idx = idx + 1) begin
                if (c_valid[idx] && !captured[idx]) begin
                    captured[idx] <= 1'b1;
                    c_flat[(idx+1)*ACC_W-1 -: ACC_W] <= c_bus[(idx+1)*ACC_W-1 -: ACC_W];
                end
            end
        end
    end

endmodule

