module pe(input clk,
            input rst,
            input[7:0] a_input,
            input[7:0] b_input,
            output[31:0] c_out
            );


for(i=0;i<=n;i++)
for(j=0;j<=m,j++)

end
ens
endmodule